i
p
pins
rotate
