cd asap7_rundir
virtuoso &

open new libr