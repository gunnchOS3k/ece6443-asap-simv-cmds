source
cd asap7_rundir
virtuoso &

